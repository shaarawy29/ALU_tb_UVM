
package my_test_pkg;
`include "test.sv"
`include "my_env.sv"
`include "my_driver.sv"
`include "my_agent.sv"
`include "my_coverage.sv"
endpackage