package my_test_pkg;
import uvm_pkg::*;
`include "my_test.sv"
`include "my_env.sv"
`include "my_driver.sv"
`include "my_agent.sv"
`include "my_coverage.sv"
`include "my_monitor.sv"
`include "my_scoreboard.sv"
`include "tx_sequence.sv"
`include "my_tx.sv"
`include "uvm_macros.svh"
`include "test_0.sv"
`include "test_transition.sv"
`include "test_1.sv"
`include "test_2.sv"
`include "test_3.sv"
`include "test_4.sv"
`include "test_5.sv"
`include "test_6.sv"
`include "test_7.sv"
`include "test_8.sv"
`include "test_9.sv"
`include "test_10.sv"
`include "test_11.sv"
`include "test_12.sv"
`include "test_13.sv"
`include "test_14.sv"
`include "test_15.sv"
endpackage