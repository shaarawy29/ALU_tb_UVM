module top_hvl;

import uvm_pkg::*;
import my_test_pkg::*;

 initial begin
 run_test();
 end

endmodule 
